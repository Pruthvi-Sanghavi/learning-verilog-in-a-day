module and_dfm(output Y, input A, B);
	assign Y = A & B;
endmodule
