module and_glm(output Y, input A, B);
	and(Y, A, B);
endmodule
